ab
aldrig
all
alla
alltid
att
av
avser
avses
bakom
bra
bredvid
de
dem
den
denna
deras
dess
det
detta
du
dä
där
efter
eftersom
efterät
ej
eller
emot
en
ett
fastän
fort
framför
från
för
genom
gott
hamske
han
hellre
hon
hos
hur
här
i
in
ingen
innan
inte
ja
jag
lite
långsamt
långt
man
med
medan
mellan
mer
mera
mindre
mot
myckett
nej
nere
ni
nu
när
nära
och
oksa
om
på
sin
skall
som
så
sådan
till
tillräckligt
tillsammans
trots
under
uppe
ut
utan
utom
vad
var
varför
vart
varthän
vem
vems
vi
vid
vilken
väl
än
ännu
är
ånyo
över
